*          Coil+ Coil- bCOM bNO bNC
.subckt DPDT  L1    L2    COM    NO   NC
S1 COM NC 10 L2 SW_NC
S2 COM NO 10 L2 SW_NO
R1 COM 0 1G
R2 NO 0 1G
R3 NC 0 1G
* R7,R8,R9,C1,D1 simulate relay operate/release delay of ~15ms
R7 L1 9 10k
R8 10 9 1meg
R9 L1 L2 1k
C1 10 L2 15nf
D1 9 L2 D
.model D D
.lib standard.dio
.model SW_NO SW(Ron=1m Roff=1G Vt=.36 Vh=.1)
.model SW_NC SW(Ron=1G Roff=1m Vt=.36 Vh=0.1)
.ends DPDT